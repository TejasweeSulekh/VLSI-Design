* Unit Inverter
.subckt inv supply Inp Output
.params widthp = 1.053u
.params widthn = 0.3161u

*Defining the parameters as a function of width
.params apd=0.18U*widthp aps=0.18U*widthp ppd=2*widthp+4*0.18U pps=2*widthp+4*0.18U
.params and=0.18U*widthn ans=0.18U*widthn pnd=2*widthn+4*0.18U pns=2*widthn+4*0.18U


* This subcircuit defines a CMOS inverter with equal n and p widths
MP1 Output Inp Supply Supply cmosp
+ L=0.18U W=widthp AD = apd AS = aps PD = ppd PS = pps
MN1 Output Inp 0 0 cmosn
+ L=0.18U W=widthn AD = and AS = ans PD = pnd PS = pns
.ends


vdd supply 0 dc 1.8

* Device under test
x3 supply Ck dutout inv

* Load Capacitor
C3 dutout 0 0.05pF

.include models-180nm

*TRANSIENT ANALYSIS with pulse inputs
VCk Ck 0 0

.dc VCk 0 1.8 0.01
.control
run
plot V(dutout)
plot deriv(dutout)
*meas tran inrise TRIG v(ck) VAL=0.18 RISE=2 TARG v(Ck) VAL=1.62 RISE=2
*meas tran infall TRIG v(ck) VAL=1.62 FALL=2 TARG v(Ck) VAL=0.18 FALL=2
*meas tran drise TRIG v(dutout) VAL=0.18 RISE=2 TARG v(dutout) VAL=1.62 RISE=2
*meas tran dfall TRIG v(dutout) VAL=1.62 FALL=2 TARG v(dutout) VAL=0.18 FALL=2
.endc
.end